module not (input in, output out);
  assign out = !in;  
endmodule